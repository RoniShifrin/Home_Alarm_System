--------------------- Title ------------------------
-- Project Name: HA_System
-- File Name: alarm_Control_TB.vhd
-- Author: Roni Shifrin
-- Ver: 1
-- Created Date: 4/12/25
----------------------------------------------------