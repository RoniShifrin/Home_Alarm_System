--------------------- Title ------------------------
-- Project Name: HA_System
-- File Name: HA_System.vhd
-- Author: Yuval Kogan
-- Ver: 1
-- Created Date: 4/12/25
----------------------------------------------------