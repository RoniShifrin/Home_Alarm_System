--------------------- Title ------------------------
-- Project Name: HA_System
-- File Name   : Alarm_controller_FSM.vhd
-- Author      : Yuval Kogan
-- Ver         : 1
-- Created Date: 04/12/25
----------------------------------------------------
